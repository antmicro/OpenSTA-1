module path_deduplication_test(
	input CLK,
	input[3:0] d,
	output[3:0] store
);
	sky130_fd_sc_hd__dfxtp_1 \store_reg[0] (
		.CLK(CLK),
		.D(d[0]),
		.Q(store[0])
	);
	
	wire store_1_inv;
	sky130_fd_sc_hd__dfxtp_1 \store_reg[1] (
		.CLK(CLK),
		.D(d[1]),
		.Q(store_1_inv)
	);
	sky130_fd_sc_hd__inv_1 _1_inv(
		.Y(store[1]),
		.A(store_1_inv)
	);

	sky130_fd_sc_hd__dfxtp_1 \store_reg[2] (
		.CLK(CLK),
		.D(d[2]),
		.Q(store[2])
	);

	sky130_fd_sc_hd__dfxtp_1 \store_reg[3] (
		.CLK(CLK),
		.D(d[3]),
		.Q(store[3])
	);
endmodule
